module ULA (
	iControl,
	iA,
	iB,
	oResult
	);

	input [4:0] iControl;
	input [31:0] iA;
	input [31:0] iB;
	output [31:0] result;
	
	always @(*)
	begin
		case (iControl)
			
		endcase
	end

endmodule